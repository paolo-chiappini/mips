
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity REGFILE is
end REGFILE;

architecture RTL of REGFILE is

begin


end RTL;

